module one_bit_comparator_structural (
    input a,
    input b,
    output greater,
    output less,
    output equal
);
    wire a_not, b_not;

    not(____); // TODO
    not(____); // TODO

    and(________); // TODO
    and(________); // TODO
    xnor(________); // TODO
endmodule
