module one_bit_comparator_behavioral (
    input a,
    input b,
    output greater,
    output less,
    output equal
);
    ____ greater = ________; // TODO
    ____ less = ________; // TODO
    ____ equal = ________; // TODO
endmodule
