module one_bit_comparator_always (
    input a,
    input b,
    output reg greater,
    output reg less,
    output reg equal
);
    always @(*) begin
        if (____) begin // TODO
            // TODO
        end else if (____) begin // TODO
            // TODO
        end else begin
            // TODO
        end
    end
endmodule
