module four_bit_comparator_always (
    input ____ a, // TODO
    input ____ b, // TODO
    output reg greater,
    output reg less,
    output reg equal
);

    always @(*) begin
        if (____) begin // TODO
            // TODO
        end else if (____) begin // TODO
            // TODO
        end else begin
            // TODO
        end
    end
endmodule
