module line_decoder (
    input [3:0] select,
    input [3:0] addr,
    output single_wire
);
    assign single_wire = ________; // TODO
endmodule
